.SUBCKT inv_1x IN OUT vm vp
*.PININFO IN:I OUT:O vm:B vp:B
MT2 OUT IN vm vm nfet W=210.0n L=60n M=1 NF=1 
MT1 OUT IN vp vp pfet W=410.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT nor3_1x A B C OUT vm vp
*.PININFO A:I B:I C:I OUT:O vm:B vp:B
MT2 OUT A vm vm nfet W=210.0n L=60n M=1 NF=1 
MT7 net010 C vp vp pfet W=810.0n L=60n M=1 NF=1 
MT3 net09 B net010 vp pfet W=810.0n L=60n M=1 NF=1 
MT1 OUT A net09 vp pfet W=810.0n L=60n M=1 NF=1 
MT8 OUT C vm vm nfet W=210.0n L=60n M=1 NF=1 
MT0 OUT B vm vm nfet W=210.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT nand2_1x A B OUT vm vp
*.PININFO A:I B:I OUT:O vm:B vp:B
MT0 net29 B vm vm nfet W=410.0n L=60n M=1 NF=1 
MT2 OUT A net29 vm nfet W=410.0n L=60n M=1 NF=1 
MT3 OUT B vp vp pfet W=410.0n L=60n M=1 NF=1 
MT1 OUT A vp vp pfet W=410.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT tgate1R_2p5u a b ng pg vm vp
*.PININFO ng:I pg:I a:B b:B vm:B vp:B
MT1 b pg a vp lvtpfet W=2.5u L=60n M=1 NF=2 
MT0 b ng a vm natnfet W=2.5u L=300n M=1 NF=2 
.ENDS

.SUBCKT R_cell3 cs gnda hmn hpn lmn lpn mo po rs vdda1p2
*.PININFO cs:I gnda:I rs:I vdda1p2:I hmn:B hpn:B lmn:B lpn:B mo:B po:B
XI1 selb sel gnda vdda1p2 / inv_1x
XI0 rs cs selb gnda vdda1p2 / nand2_1x
RR2 hpn lpn r=60.08182 
RR0 lmn hmn r=60.08182 
XI3 lmn mo sel selb gnda vdda1p2 / tgate1R_2p5u
XI2 lpn po sel selb gnda vdda1p2 / tgate1R_2p5u
.ENDS

.SUBCKT R_array2 B<5> B<4> B<3> B<2> B<1> B<0> gnda im ip mo po vcm vdda1p2
*.PININFO B<5>:I B<4>:I B<3>:I B<2>:I B<1>:I B<0>:I gnda:I im:I ip:I vcm:I 
*.PININFO vdda1p2:I mo:O po:O
XI85 B<0> Bb<0> gnda vdda1p2 / inv_1x
XI84 B<1> Bb<1> gnda vdda1p2 / inv_1x
XI83 B<2> Bb<2> gnda vdda1p2 / inv_1x
XI82 B<3> Bb<3> gnda vdda1p2 / inv_1x
XI81 B<4> Bb<4> gnda vdda1p2 / inv_1x
XI80 B<5> Bb<5> gnda vdda1p2 / inv_1x
XI79 Bb<5> Bb<4> Bb<3> net11 gnda vdda1p2 / nor3_1x
XI78 Bb<5> Bb<4> B<3> net12 gnda vdda1p2 / nor3_1x
XI77 Bb<5> B<4> Bb<3> net13 gnda vdda1p2 / nor3_1x
XI76 Bb<5> B<4> B<3> net14 gnda vdda1p2 / nor3_1x
XI75 B<5> Bb<4> Bb<3> net15 gnda vdda1p2 / nor3_1x
XI74 B<5> Bb<4> B<3> net16 gnda vdda1p2 / nor3_1x
XI73 B<5> B<4> Bb<3> net17 gnda vdda1p2 / nor3_1x
XI72 B<5> B<4> B<3> net18 gnda vdda1p2 / nor3_1x
XI71 Bb<2> Bb<1> Bb<0> net39 gnda vdda1p2 / nor3_1x
XI70 Bb<2> Bb<1> B<0> net36 gnda vdda1p2 / nor3_1x
XI69 Bb<2> B<1> Bb<0> net33 gnda vdda1p2 / nor3_1x
XI68 Bb<2> B<1> B<0> net30 gnda vdda1p2 / nor3_1x
XI67 B<2> Bb<1> Bb<0> net27 gnda vdda1p2 / nor3_1x
XI66 B<2> Bb<1> B<0> net24 gnda vdda1p2 / nor3_1x
XI65 B<2> B<1> Bb<0> net21 gnda vdda1p2 / nor3_1x
XI64 B<2> B<1> B<0> net10 gnda vdda1p2 / nor3_1x
XI63 net10 gnda net297 net298 net82 net74 mo po net14 vdda1p2 / R_cell3
XI62 net10 gnda net281 net282 net84 net76 mo po net12 vdda1p2 / R_cell3
XI61 net10 gnda net255 net256 net85 net77 mo po net11 vdda1p2 / R_cell3
XI60 net30 gnda net247 net248 net249 net250 mo po net11 vdda1p2 / R_cell3
XI59 net36 gnda net243 net244 net245 net246 mo po net11 vdda1p2 / R_cell3
XI58 net39 gnda im ip net243 net244 mo po net11 vdda1p2 / R_cell3
XI57 net33 gnda net245 net246 net247 net248 mo po net11 vdda1p2 / R_cell3
XI56 net24 gnda net251 net252 net253 net254 mo po net11 vdda1p2 / R_cell3
XI55 net27 gnda net249 net250 net251 net252 mo po net11 vdda1p2 / R_cell3
XI54 net21 gnda net253 net254 net255 net256 mo po net11 vdda1p2 / R_cell3
XI53 net30 gnda net265 net266 net269 net270 mo po net12 vdda1p2 / R_cell3
XI52 net36 gnda net257 net258 net261 net262 mo po net12 vdda1p2 / R_cell3
XI51 net39 gnda net85 net77 net257 net258 mo po net12 vdda1p2 / R_cell3
XI50 net33 gnda net261 net262 net265 net266 mo po net12 vdda1p2 / R_cell3
XI49 net24 gnda net273 net274 net277 net278 mo po net12 vdda1p2 / R_cell3
XI48 net27 gnda net269 net270 net273 net274 mo po net12 vdda1p2 / R_cell3
XI47 net21 gnda net277 net278 net281 net282 mo po net12 vdda1p2 / R_cell3
XI46 net10 gnda net283 net284 net83 net75 mo po net13 vdda1p2 / R_cell3
XI45 net30 gnda net267 net268 net271 net272 mo po net13 vdda1p2 / R_cell3
XI44 net36 gnda net259 net260 net263 net264 mo po net13 vdda1p2 / R_cell3
XI43 net39 gnda net84 net76 net259 net260 mo po net13 vdda1p2 / R_cell3
XI42 net33 gnda net263 net264 net267 net268 mo po net13 vdda1p2 / R_cell3
XI41 net24 gnda net275 net276 net279 net280 mo po net13 vdda1p2 / R_cell3
XI40 net27 gnda net271 net272 net275 net276 mo po net13 vdda1p2 / R_cell3
XI39 net21 gnda net279 net280 net283 net284 mo po net13 vdda1p2 / R_cell3
XI38 net30 gnda net289 net290 net291 net292 mo po net14 vdda1p2 / R_cell3
XI37 net36 gnda net285 net286 net287 net288 mo po net14 vdda1p2 / R_cell3
XI36 net39 gnda net83 net75 net285 net286 mo po net14 vdda1p2 / R_cell3
XI35 net33 gnda net287 net288 net289 net290 mo po net14 vdda1p2 / R_cell3
XI34 net24 gnda net293 net294 net295 net296 mo po net14 vdda1p2 / R_cell3
XI33 net27 gnda net291 net292 net293 net294 mo po net14 vdda1p2 / R_cell3
XI32 net21 gnda net295 net296 net297 net298 mo po net14 vdda1p2 / R_cell3
XI31 net10 gnda net325 net326 net80 net72 mo po net16 vdda1p2 / R_cell3
XI30 net10 gnda net311 net312 net81 net73 mo po net15 vdda1p2 / R_cell3
XI29 net30 gnda net303 net304 net305 net306 mo po net15 vdda1p2 / R_cell3
XI28 net36 gnda net299 net300 net301 net302 mo po net15 vdda1p2 / R_cell3
XI27 net39 gnda net82 net74 net299 net300 mo po net15 vdda1p2 / R_cell3
XI26 net33 gnda net301 net302 net303 net304 mo po net15 vdda1p2 / R_cell3
XI25 net24 gnda net307 net308 net309 net310 mo po net15 vdda1p2 / R_cell3
XI24 net27 gnda net305 net306 net307 net308 mo po net15 vdda1p2 / R_cell3
XI23 net21 gnda net309 net310 net311 net312 mo po net15 vdda1p2 / R_cell3
XI22 net30 gnda net317 net318 net319 net320 mo po net16 vdda1p2 / R_cell3
XI21 net36 gnda net313 net314 net315 net316 mo po net16 vdda1p2 / R_cell3
XI20 net39 gnda net81 net73 net313 net314 mo po net16 vdda1p2 / R_cell3
XI19 net33 gnda net315 net316 net317 net318 mo po net16 vdda1p2 / R_cell3
XI18 net24 gnda net321 net322 net323 net324 mo po net16 vdda1p2 / R_cell3
XI17 net27 gnda net319 net320 net321 net322 mo po net16 vdda1p2 / R_cell3
XI16 net21 gnda net323 net324 net325 net326 mo po net16 vdda1p2 / R_cell3
XI15 net10 gnda net339 net340 net79 net71 mo po net17 vdda1p2 / R_cell3
XI14 net30 gnda net331 net332 net333 net334 mo po net17 vdda1p2 / R_cell3
XI13 net36 gnda net327 net328 net329 net330 mo po net17 vdda1p2 / R_cell3
XI12 net39 gnda net80 net72 net327 net328 mo po net17 vdda1p2 / R_cell3
XI11 net33 gnda net329 net330 net331 net332 mo po net17 vdda1p2 / R_cell3
XI10 net24 gnda net335 net336 net337 net338 mo po net17 vdda1p2 / R_cell3
XI9 net27 gnda net333 net334 net335 net336 mo po net17 vdda1p2 / R_cell3
XI8 net21 gnda net337 net338 net339 net340 mo po net17 vdda1p2 / R_cell3
XI7 net30 gnda net345 net346 net347 net348 mo po net18 vdda1p2 / R_cell3
XI6 net36 gnda net341 net342 net343 net344 mo po net18 vdda1p2 / R_cell3
XI5 net39 gnda net79 net71 net341 net342 mo po net18 vdda1p2 / R_cell3
XI4 net33 gnda net343 net344 net345 net346 mo po net18 vdda1p2 / R_cell3
XI3 net24 gnda net349 net350 net351 net352 mo po net18 vdda1p2 / R_cell3
XI2 net27 gnda net347 net348 net349 net350 mo po net18 vdda1p2 / R_cell3
XI1 net21 gnda net351 net352 net353 net354 mo po net18 vdda1p2 / R_cell3
XI0 net10 gnda net353 net354 vcm vcm mo po net18 vdda1p2 / R_cell3
.ENDS

.SUBCKT tgate1R_p5u a b ng pg vm vp
*.PININFO ng:I pg:I a:B b:B vm:B vp:B
MT1 b pg a vp lvtpfet W=500n L=60n M=1 NF=1 
MT0 b ng a vm natnfet W=500n L=300n M=1 NF=1 
.ENDS

.SUBCKT cap_cell_dummy2 vcm vm vp
*.PININFO vcm:I vm:I vp:I
XI11 sel sb posb vm vp / nand2_1x
XI8 sel vm negb vm vp / nand2_1x
XI5 vm net026 sel vm vp / nand2_1x
XI0 vm vm net026 vm vp / nand2_1x
MT1 vcm selb net19 vm nfet W=210.0n L=60n M=1 NF=1 
MT0 net21 selb vcm vm nfet W=210.0n L=60n M=1 NF=1 
CC1 vm net19 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
CC0 vm net21 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
XI12 vm sb vm vp / inv_1x
XI10 posb pos vm vp / inv_1x
XI9 negb neg vm vp / inv_1x
XI2 sel selb vm vp / inv_1x
XI7 vm net19 neg negb vm vp / tgate1R_p5u
XI6 vm net21 neg negb vm vp / tgate1R_p5u
XI4 vm net19 pos posb vm vp / tgate1R_p5u
XI3 vm net21 pos posb vm vp / tgate1R_p5u
.ENDS

.SUBCKT tgateL1p5R a b ng pg vm vp
*.PININFO ng:I pg:I a:B b:B vm:B vp:B
MT1 b pg a vp lvtpfet W=137.5u L=60n M=1 NF=22 
MT0 b ng a vm natnfet W=124.74u L=300n M=1 NF=22 
.ENDS

.SUBCKT cap_cell2 am ap c im ip nrb r s vcm vm vp
*.PININFO c:I im:I ip:I nrb:I r:I s:I vcm:I vm:I vp:I am:B ap:B
XI12 s sb vm vp / inv_1x
XI10 posb pos vm vp / inv_1x
XI9 negb neg vm vp / inv_1x
XI2 sel selb vm vp / inv_1x
XI11 sel sb posb vm vp / nand2_1x
XI8 sel s negb vm vp / nand2_1x
XI5 nrb net026 sel vm vp / nand2_1x
XI0 r c net026 vm vp / nand2_1x
CC1 ap net19 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
CC0 am net21 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
XI7 ip net19 neg negb vm vp / tgate1R_p5u
XI6 im net21 neg negb vm vp / tgate1R_p5u
XI4 im net19 pos posb vm vp / tgate1R_p5u
XI16 vcm net21 selb sel vm vp / tgate1R_p5u
XI17 vcm net19 selb sel vm vp / tgate1R_p5u
XI3 ip net21 pos posb vm vp / tgate1R_p5u
.ENDS

.SUBCKT cap_cell_tr am ap im ip p1 p2 s vcm vm vp
*.PININFO im:I ip:I p1:I p2:I s:I vcm:I vm:I vp:I am:B ap:B
XI11 p2 sb posb vm vp / nand2_1x
XI8 p2 s negb vm vp / nand2_1x
XI12 s sb vm vp / inv_1x
XI10 posb pos vm vp / inv_1x
XI9 negb neg vm vp / inv_1x
XI17 p1 p1b vm vp / inv_1x
CC1 ap net19 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
CC0 am net21 $[vncap] $SUB=vm w=6.9u l=7u botlev=2 toplev=5 setind=-1.0
XI7 ip net19 neg negb vm vp / tgate1R_p5u
XI6 im net21 neg negb vm vp / tgate1R_p5u
XI4 im net19 pos posb vm vp / tgate1R_p5u
XI16 vcm net21 p1 p1b vm vp / tgate1R_p5u
XI3 ip net21 pos posb vm vp / tgate1R_p5u
XI19 vcm net19 p1 p1b vm vp / tgate1R_p5u
.ENDS

.SUBCKT nor2_1x A B OUT vm vp
*.PININFO A:I B:I OUT:O vm:B vp:B
MT0 OUT B vm vm nfet W=210.0n L=60n M=1 NF=1 
MT2 OUT A vm vm nfet W=210.0n L=60n M=1 NF=1 
MT3 net09 A vp vp pfet W=810.0n L=60n M=1 NF=1 
MT1 OUT B net09 vp pfet W=810.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT inv_32x IN OUT vm vp
*.PININFO IN:I OUT:O vm:B vp:B
MT2 OUT IN vm vm nfet W=6.56u L=60n M=1 NF=16 
MT1 OUT IN vp vp pfet W=12.96u L=60n M=1 NF=16 
.ENDS

.SUBCKT nand3_1x A B C OUT vm vp
*.PININFO A:I B:I C:I OUT:O vm:B vp:B
MT5 net27 C vm vm nfet W=410.0n L=60n M=1 NF=1 
MT0 net29 B net27 vm nfet W=410.0n L=60n M=1 NF=1 
MT2 OUT A net29 vm nfet W=410.0n L=60n M=1 NF=1 
MT4 OUT C vp vp pfet W=410.0n L=60n M=1 NF=1 
MT3 OUT B vp vp pfet W=410.0n L=60n M=1 NF=1 
MT1 OUT A vp vp pfet W=410.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT cap_array5 B<12> B<11> B<10> B<9> B<8> B<7> B<6> BC Ho Sa am ap gnda 
+ im ip lam lap refm refp vcm vdda1p2
*.PININFO B<12>:I B<11>:I B<10>:I B<9>:I B<8>:I B<7>:I B<6>:I BC:I Ho:I Sa:I 
*.PININFO gnda:I im:I ip:I lam:I lap:I refm:I refp:I vcm:I vdda1p2:I am:B ap:B
XI179 net0402 SaHo gnda vdda1p2 / inv_1x
XI102 B<6> Bb<6> gnda vdda1p2 / inv_1x
XI101 B<7> Bb<7> gnda vdda1p2 / inv_1x
XI100 B<9> Bb<9> gnda vdda1p2 / inv_1x
XI99 B<8> Bb<8> gnda vdda1p2 / inv_1x
XI98 B<10> Bb<10> gnda vdda1p2 / inv_1x
XI97 B<11> Bb<11> gnda vdda1p2 / inv_1x
XI165 net16 net038 gnda vdda1p2 / inv_1x
XI166 net6 net033 gnda vdda1p2 / inv_1x
XI175 Sab net0396 gnda vdda1p2 / inv_1x
XI162 net239 net034 gnda vdda1p2 / inv_1x
XI163 net10 net035 gnda vdda1p2 / inv_1x
XI164 net14 net037 gnda vdda1p2 / inv_1x
XI167 net20 net039 gnda vdda1p2 / inv_1x
XI95 Bb<6> Bb<7> Bb<8> net0266 gnda vdda1p2 / nor3_1x
XI79 Bb<9> Bb<10> Bb<11> net20 gnda vdda1p2 / nor3_1x
XI168<1> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<2> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<3> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<4> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<5> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<6> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<7> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<8> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<9> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<10> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<11> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<12> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<13> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<14> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<15> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<16> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<17> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<18> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<19> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<20> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<21> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<22> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<23> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<24> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<25> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<26> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<27> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<28> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<29> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<30> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<31> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<32> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<33> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<34> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<35> vcm gnda vdda1p2 / cap_cell_dummy2
XI168<36> vcm gnda vdda1p2 / cap_cell_dummy2
XI174 am vcm Sa Sab gnda vdda1p2 / tgateL1p5R
XI173 ap vcm Sa Sab gnda vdda1p2 / tgateL1p5R
XI170 cip refp BC BCb gnda vdda1p2 / tgateL1p5R
XI151 cip ip Sai Saib gnda vdda1p2 / tgateL1p5R
XI171 cim refm BC BCb gnda vdda1p2 / tgateL1p5R
XI153 cim im Sai Saib gnda vdda1p2 / tgateL1p5R
XI63 am ap net4 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI62 am ap net4 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI61 am ap net4 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI60 am ap net0268 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI59 am ap net0266 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI57 am ap net0267 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI56 am ap net0271 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI55 am ap B<8> cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI54 am ap net25 cim cip vdda1p2 net20 B<12> vcm gnda vdda1p2 / cap_cell2
XI53 am ap net0268 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI52 am ap net0266 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI51 am ap gnda cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI50 am ap net0267 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI49 am ap net0271 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI48 am ap B<8> cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI47 am ap net25 cim cip net039 net16 B<12> vcm gnda vdda1p2 / cap_cell2
XI46 am ap net4 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI45 am ap net0268 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI44 am ap net0266 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI43 am ap gnda cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI42 am ap net0267 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI41 am ap net0271 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI40 am ap B<8> cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI39 am ap net25 cim cip net038 net14 B<12> vcm gnda vdda1p2 / cap_cell2
XI38 am ap net0268 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI37 am ap net0266 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI36 am ap gnda cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI35 am ap net0267 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI34 am ap net0271 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI33 am ap B<8> cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI32 am ap net25 cim cip net037 B<11> B<12> vcm gnda vdda1p2 / cap_cell2
XI31 am ap net4 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI30 am ap net4 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI29 am ap net0268 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI28 am ap net0266 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI27 am ap gnda cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI26 am ap net0267 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI25 am ap net0271 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI24 am ap B<8> cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI23 am ap net25 cim cip Bb<11> net10 B<12> vcm gnda vdda1p2 / cap_cell2
XI22 am ap net0268 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI21 am ap net0266 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI20 am ap gnda cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI19 am ap net0267 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI18 am ap net0271 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI17 am ap B<8> cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI16 am ap net25 cim cip net035 net239 B<12> vcm gnda vdda1p2 / cap_cell2
XI15 am ap net4 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI14 am ap net0268 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI13 am ap net0266 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI12 am ap gnda cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI11 am ap net0267 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI10 am ap net0271 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI9 am ap B<8> cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI8 am ap net25 cim cip net034 net6 B<12> vcm gnda vdda1p2 / cap_cell2
XI7 am ap net0268 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI6 am ap net0266 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI5 am ap gnda cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI4 am ap net0267 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI3 am ap net0271 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI2 am ap B<8> cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI1 am ap net25 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI0 am ap net4 cim cip net033 vdda1p2 B<12> vcm gnda vdda1p2 / cap_cell2
XI58 am ap lam lap SaHo BC B<12> vcm gnda vdda1p2 / cap_cell_tr
XI178 Ho net0396 net0402 gnda vdda1p2 / nor2_1x
XI94 Bb<8> Bb<7> net0267 gnda vdda1p2 / nor2_1x
XI93 B<7> B<6> net0269 gnda vdda1p2 / nor2_1x
XI92 Bb<8> net0269 net0268 gnda vdda1p2 / nor2_1x
XI78 Bb<11> Bb<10> net16 gnda vdda1p2 / nor2_1x
XI77 B<10> B<9> net227 gnda vdda1p2 / nor2_1x
XI76 Bb<11> net227 net14 gnda vdda1p2 / nor2_1x
XI91 B<7> B<6> net0270 gnda vdda1p2 / nand2_1x
XI90 Bb<8> net0270 net0271 gnda vdda1p2 / nand2_1x
XI89 Bb<8> Bb<7> net25 gnda vdda1p2 / nand2_1x
XI75 Bb<11> Bb<10> net239 gnda vdda1p2 / nand2_1x
XI74 B<10> B<9> net238 gnda vdda1p2 / nand2_1x
XI73 Bb<11> net238 net10 gnda vdda1p2 / nand2_1x
XI172 BC BCb gnda vdda1p2 / inv_32x
XI177 Saib Sai gnda vdda1p2 / inv_32x
XI176 net0396 Saib gnda vdda1p2 / inv_32x
XI156 Sa Sab gnda vdda1p2 / inv_32x
XI88 Bb<8> Bb<7> Bb<6> net4 gnda vdda1p2 / nand3_1x
XI72 Bb<11> Bb<10> Bb<9> net6 gnda vdda1p2 / nand3_1x
.ENDS

.SUBCKT DAC_array B<12> B<11> B<10> B<9> B<8> B<7> B<6> B<5> B<4> B<3> B<2> 
+ B<1> B<0> BC Ho Sa am ap gnda im ip refm refp vcm vdda1p2
*.PININFO B<12>:I B<11>:I B<10>:I B<9>:I B<8>:I B<7>:I B<6>:I B<5>:I B<4>:I 
*.PININFO B<3>:I B<2>:I B<1>:I B<0>:I BC:I Ho:I Sa:I gnda:I im:I ip:I refm:I 
*.PININFO refp:I vcm:I vdda1p2:I am:B ap:B
XI2 B<5> B<4> B<3> B<2> B<1> B<0> gnda refm refp lam lap vcm vdda1p2 / R_array2
XI1 B<12> B<11> B<10> B<9> B<8> B<7> B<6> BC Ho Sa am ap gnda im ip lam lap 
+ refm refp vcm vdda1p2 / cap_array5
.ENDS

.SUBCKT inv_8x IN OUT vm vp
*.PININFO IN:I OUT:O vm:B vp:B
MT2 OUT IN vm vm nfet W=1.64u L=60n M=1 NF=4 
MT1 OUT IN vp vp pfet W=3.24u L=60n M=1 NF=4 
.ENDS

.SUBCKT sarc B Cob Cp Ho Npb S ckb gnd vdd1p2
*.PININFO Cob:I Cp:I Ho:I Npb:I S:I ckb:I B:O gnd:B vdd1p2:B
XI3 net15 B gnd vdd1p2 / inv_8x
XI2 Cob ckb Npb net21 gnd vdd1p2 / nor3_1x
XI1 net21 Ho net15 net012 gnd vdd1p2 / nor3_1x
XI0 Cp net012 S net15 gnd vdd1p2 / nor3_1x
.ENDS

.SUBCKT tgate0 a b ng pg vm vp
*.PININFO ng:I pg:I a:B b:B vm:B vp:B
MT0 b ng a vm nfet W=210.0n L=60n M=1 NF=1 
MT1 b pg a vp pfet W=410.0n L=60n M=1 NF=1 
.ENDS

.SUBCKT inv_4x IN OUT vm vp
*.PININFO IN:I OUT:O vm:B vp:B
MT2 OUT IN vm vm nfet W=820.0n L=60n M=1 NF=2 
MT1 OUT IN vp vp pfet W=1.62u L=60n M=1 NF=2 
.ENDS

.SUBCKT dffr CK D Q Qb RN vm vp
*.PININFO CK:I D:I RN:I vm:I vp:I Q:O Qb:O
XI6 net16 net14 clk clkb vm vp / tgate0
XI5 net52 net16 clkb clk vm vp / tgate0
XI4 net53 net13 clk clkb vm vp / tgate0
XI1 net54 net13 clkb clk vm vp / tgate0
XI12 clkb clk vm vp / inv_1x
XI11 CK clkb vm vp / inv_1x
XI10 Q Qb vm vp / inv_1x
XI9 net17 Q vm vp / inv_1x
XI8 net17 net52 vm vp / inv_1x
XI2 net13 net14 vm vp / inv_1x
XI0 D net54 vm vp / inv_1x
XI7 net16 RN net17 vm vp / nand2_1x
XI3 RN net14 net53 vm vp / nand2_1x
.ENDS

.SUBCKT dffs CK D Q Qb SN vm vp
*.PININFO CK:I D:I SN:I vm:I vp:I Q:O Qb:O
XI12 clkb clk vm vp / inv_1x
XI11 CK clkb vm vp / inv_1x
XI10 Q Qb vm vp / inv_1x
XI9 net17 Q vm vp / inv_1x
XI7 net16 net17 vm vp / inv_1x
XI3 net14 net53 vm vp / inv_1x
XI0 D net54 vm vp / inv_1x
XI8 net17 SN net52 vm vp / nand2_1x
XI2 SN net13 net14 vm vp / nand2_1x
XI6 net16 net52 clkb clk vm vp / tgate0
XI5 net14 net16 clk clkb vm vp / tgate0
XI4 net53 net13 clk clkb vm vp / tgate0
XI1 net54 net13 clkb clk vm vp / tgate0
.ENDS

.SUBCKT Shf_line Q<13> Q<12> Q<11> Q<10> Q<9> Q<8> Q<7> Q<6> Q<5> Q<4> Q<3> 
+ Q<2> Q<1> Q<0> Qb<13> Qb<12> Qb<11> Qb<10> Qb<9> Qb<8> Qb<7> Qb<6> Qb<5> 
+ Qb<4> Qb<3> Qb<2> Qb<1> Qb<0> RN ck ckbbf ckl cko gnd vdd1p2
*.PININFO RN:I ck:I gnd:I vdd1p2:I Q<13>:O Q<12>:O Q<11>:O Q<10>:O Q<9>:O 
*.PININFO Q<8>:O Q<7>:O Q<6>:O Q<5>:O Q<4>:O Q<3>:O Q<2>:O Q<1>:O Q<0>:O 
*.PININFO Qb<13>:O Qb<12>:O Qb<11>:O Qb<10>:O Qb<9>:O Qb<8>:O Qb<7>:O Qb<6>:O 
*.PININFO Qb<5>:O Qb<4>:O Qb<3>:O Qb<2>:O Qb<1>:O Qb<0>:O ckbbf:O ckl:O cko:O
XI13 net07 net18 Q<13> Qb<13> net8 gnd vdd1p2 / dffr
XI12 net07 Q<13> Q<12> Qb<12> net8 gnd vdd1p2 / dffr
XI11 net07 Q<12> Q<11> Qb<11> net8 gnd vdd1p2 / dffr
XI10 net07 Q<11> Q<10> Qb<10> net8 gnd vdd1p2 / dffr
XI9 net07 Q<10> Q<9> Qb<9> net8 gnd vdd1p2 / dffr
XI8 net07 Q<9> Q<8> Qb<8> net8 gnd vdd1p2 / dffr
XI7 net07 Q<8> Q<7> Qb<7> net8 gnd vdd1p2 / dffr
XI6 net07 Q<7> Q<6> Qb<6> net8 gnd vdd1p2 / dffr
XI5 net07 Q<6> Q<5> Qb<5> net8 gnd vdd1p2 / dffr
XI4 net07 Q<5> Q<4> Qb<4> net8 gnd vdd1p2 / dffr
XI3 net07 Q<4> Q<3> Qb<3> net8 gnd vdd1p2 / dffr
XI2 net07 Q<3> Q<2> Qb<2> net8 gnd vdd1p2 / dffr
XI1 net07 Q<2> Q<1> Qb<1> net8 gnd vdd1p2 / dffr
XI31 net026 net031 gnd vdd1p2 / inv_1x
XI30 net020 net026 gnd vdd1p2 / inv_1x
XI29 net023 net022 gnd vdd1p2 / inv_1x
XI28 net031 net023 gnd vdd1p2 / inv_1x
XI26 net023 cko gnd vdd1p2 / inv_1x
XI25 net019 net020 gnd vdd1p2 / inv_1x
XI24 net07 net019 gnd vdd1p2 / inv_1x
XI18 net19 net18 gnd vdd1p2 / inv_1x
XI17 Q<0> net19 gnd vdd1p2 / inv_1x
XI27 net022 ckbbf gnd vdd1p2 / inv_4x
XI21 RN net20 gnd vdd1p2 / inv_4x
XI19 ck net21 gnd vdd1p2 / inv_4x
XI22 net20 net8 gnd vdd1p2 / inv_32x
XI20 net21 net07 gnd vdd1p2 / inv_32x
XI0 net07 Q<1> Q<0> Qb<0> net8 gnd vdd1p2 / dffs
XI33 net032 Q<13> net038 gnd vdd1p2 / nor2_1x
XI32 Qb<13> net21 net032 gnd vdd1p2 / nor2_1x
XI34 net038 ckl gnd vdd1p2 / inv_8x
.ENDS

.SUBCKT sarlogic2 ADCo BC Co Cob D<11> D<10> D<9> D<8> D<7> D<6> D<5> D<4> 
+ D<3> D<2> D<1> D<0> Ho PO<11> PO<10> PO<9> PO<8> PO<7> PO<6> PO<5> PO<4> 
+ PO<3> PO<2> PO<1> PO<0> RN Sa ck gnd lat vdd1p2 vddp
*.PININFO Co:I Cob:I RN:I ck:I ADCo:O BC:O D<11>:O D<10>:O D<9>:O D<8>:O 
*.PININFO D<7>:O D<6>:O D<5>:O D<4>:O D<3>:O D<2>:O D<1>:O D<0>:O Ho:O 
*.PININFO PO<11>:O PO<10>:O PO<9>:O PO<8>:O PO<7>:O PO<6>:O PO<5>:O PO<4>:O 
*.PININFO PO<3>:O PO<2>:O PO<1>:O PO<0>:O Sa:O lat:O gnd:B vdd1p2:B vddp:B
XI5 Q<10> net17 net11 gnd vdd1p2 / nor2_1x
XI2 Q<11> net13 net015 gnd vdd1p2 / nor2_1x
XI1 Q<13> net015 net13 gnd vdd1p2 / nor2_1x
XI23<11> net063<0> PO<11> gnd vddp / inv_32x
XI23<10> net063<1> PO<10> gnd vddp / inv_32x
XI23<9> net063<2> PO<9> gnd vddp / inv_32x
XI23<8> net063<3> PO<8> gnd vddp / inv_32x
XI23<7> net063<4> PO<7> gnd vddp / inv_32x
XI23<6> net063<5> PO<6> gnd vddp / inv_32x
XI23<5> net063<6> PO<5> gnd vddp / inv_32x
XI23<4> net063<7> PO<4> gnd vddp / inv_32x
XI23<3> net063<8> PO<3> gnd vddp / inv_32x
XI23<2> net063<9> PO<2> gnd vddp / inv_32x
XI23<1> net063<10> PO<1> gnd vddp / inv_32x
XI23<0> net063<11> PO<0> gnd vddp / inv_32x
XI8 net074 BC gnd vdd1p2 / inv_32x
XI4 net41 Ho gnd vdd1p2 / inv_32x
XI172 net13 Sa gnd vdd1p2 / inv_32x
XI28 Qb<11> net17 net074 gnd vdd1p2 / nand2_1x
XI3 Q<11> net029 net41 gnd vdd1p2 / nand2_1x
XI6 Q<13> net11 net40 net17 gnd vdd1p2 / nor3_1x
XI27 D<11> Db<11> gnd vdd1p2 / inv_1x
XI13 Q<0> net041 gnd vdd1p2 / inv_1x
XI14 Sa net029 gnd vdd1p2 / inv_1x
XI7 RN net40 gnd vdd1p2 / inv_1x
XI9<10> D<10> ACo Q<10> Ho Qb<9> Sa lat gnd vdd1p2 / sarc
XI9<9> D<9> ACo Q<9> Ho Qb<8> Sa lat gnd vdd1p2 / sarc
XI9<8> D<8> ACo Q<8> Ho Qb<7> Sa lat gnd vdd1p2 / sarc
XI9<7> D<7> ACo Q<7> Ho Qb<6> Sa lat gnd vdd1p2 / sarc
XI9<6> D<6> ACo Q<6> Ho Qb<5> Sa lat gnd vdd1p2 / sarc
XI9<5> D<5> ACo Q<5> Ho Qb<4> Sa lat gnd vdd1p2 / sarc
XI9<4> D<4> ACo Q<4> Ho Qb<3> Sa lat gnd vdd1p2 / sarc
XI9<3> D<3> ACo Q<3> Ho Qb<2> Sa lat gnd vdd1p2 / sarc
XI9<2> D<2> ACo Q<2> Ho Qb<1> Sa lat gnd vdd1p2 / sarc
XI9<1> D<1> ACo Q<1> Ho Qb<0> Sa lat gnd vdd1p2 / sarc
XI15 D<11> Cob Q<11> gnd Qb<10> Sa lat gnd vdd1p2 / sarc
XI25 Co net082 D<11> Db<11> gnd vdd1p2 / tgate0
XI24 Cob net082 Db<11> D<11> gnd vdd1p2 / tgate0
XI26 net082 ACo gnd vdd1p2 / inv_4x
XI12 net041 D<0> gnd vdd1p2 / inv_4x
XI22<11> ckl D<11> net069<0> net063<0> RN gnd vdd1p2 / dffr
XI22<10> ckl D<10> net069<1> net063<1> RN gnd vdd1p2 / dffr
XI22<9> ckl D<9> net069<2> net063<2> RN gnd vdd1p2 / dffr
XI22<8> ckl D<8> net069<3> net063<3> RN gnd vdd1p2 / dffr
XI22<7> ckl D<7> net069<4> net063<4> RN gnd vdd1p2 / dffr
XI22<6> ckl D<6> net069<5> net063<5> RN gnd vdd1p2 / dffr
XI22<5> ckl D<5> net069<6> net063<6> RN gnd vdd1p2 / dffr
XI22<4> ckl D<4> net069<7> net063<7> RN gnd vdd1p2 / dffr
XI22<3> ckl D<3> net069<8> net063<8> RN gnd vdd1p2 / dffr
XI22<2> ckl D<2> net069<9> net063<9> RN gnd vdd1p2 / dffr
XI22<1> ckl D<1> net069<10> net063<10> RN gnd vdd1p2 / dffr
XI22<0> ckl ACo net069<11> net063<11> RN gnd vdd1p2 / dffr
XI19 cko Co ADCo net055 RN gnd vdd1p2 / dffr
XI0 Q<13> Q<12> Q<11> Q<10> Q<9> Q<8> Q<7> Q<6> Q<5> Q<4> Q<3> Q<2> Q<1> Q<0> 
+ Qb<13> Qb<12> Qb<11> Qb<10> Qb<9> Qb<8> Qb<7> Qb<6> Qb<5> Qb<4> Qb<3> Qb<2> 
+ Qb<1> Qb<0> RN ck lat ckl cko gnd vdd1p2 / Shf_line
.ENDS

.SUBCKT comp2 gnda ib im ip lat om on op vdda1p2
*.PININFO gnda:I ib:I im:I ip:I lat:I on:I vdda1p2:I om:O op:O
MT29 net0138 on gnda gnda nfet W=10u L=60n M=1 NF=2 
MT19 net035 lat net0138 gnda nfet W=6u L=60n M=1 NF=2 
RR1 o1m net49 r=12.75K 
RR0 net49 o1p r=12.75K 
MT4 o1p net49 vdda1p2 vdda1p2 pfet W=40u L=500n M=1 NF=8 
MT3 o1m net49 vdda1p2 vdda1p2 pfet W=40u L=500n M=1 NF=8 
MT27 vdda1p2 o1p o1pbf gnda natnfet W=20u L=300n M=1 NF=4 
MT24 vdda1p2 o1m o1mbf gnda natnfet W=20u L=300n M=1 NF=4 
MT2 o1m ip net47 gnda natnfet W=15.0u L=300n M=1 NF=3 
MT1 o1p im net47 gnda natnfet W=15.0u L=300n M=1 NF=3 
MT16 rgm rgp net035 gnda nfet W=10u L=600n M=1 NF=2 
MT15 rgp rgm net035 gnda nfet W=10u L=600n M=1 NF=2 
MT17 rgm o1pbf vdda1p2 vdda1p2 lvtpfet W=9u L=600n M=1 NF=3 
MT14 rgp o1mbf vdda1p2 vdda1p2 lvtpfet W=9u L=600n M=1 NF=3 
MT30 ib onb vbn vdda1p2 pfet W=5u L=60n M=1 NF=1 
MT54 gnda onb vbn gnda nfet W=5u L=60n M=1 NF=1 
MT26 o1pbf vbn gnda gnda nfet W=10u L=500n M=6 NF=2 
MT25 o1mbf vbn gnda gnda nfet W=10u L=500n M=6 NF=2 
MT20 vbn vbn gnda gnda nfet W=10u L=500n M=1 NF=2 
MT0 net47 vbn gnda gnda nfet W=10u L=500n M=20 NF=2 
XI1 rgp op om gnda vdda1p2 / nand2_1x
XI0 rgm om op gnda vdda1p2 / nand2_1x
MT21 rgp lat vdda1p2 vdda1p2 lvtpfet W=500n L=60n M=1 NF=1 
MT18 rgm lat vdda1p2 vdda1p2 lvtpfet W=500n L=60n M=1 NF=1 
MT31 gnda vbn gnda gnda nfet W=85.0u L=5u M=1 NF=17 
XI17 on onb gnda vdda1p2 / inv_1x
.ENDS

.SUBCKT ADC12b ADCo Ho PO<11> PO<10> PO<9> PO<8> PO<7> PO<6> PO<5> PO<4> PO<3> 
+ PO<2> PO<1> PO<0> RN ck gnd ib im ip on refm refp sync vcm vdd1p2 vdda1p2 
+ vddp
*.PININFO RN:I ck:I ib:I im:I ip:I on:I refm:I refp:I vcm:I ADCo:O Ho:O 
*.PININFO PO<11>:O PO<10>:O PO<9>:O PO<8>:O PO<7>:O PO<6>:O PO<5>:O PO<4>:O 
*.PININFO PO<3>:O PO<2>:O PO<1>:O PO<0>:O sync:O gnd:B vdd1p2:B vdda1p2:B 
*.PININFO vddp:B
XI1 D<11> D<10> D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> D<0> gnd BC Ho Sa 
+ am ap gnd im ip refm refp vcm vdda1p2 / DAC_array
XI3 BC net44 gnd vddp / inv_1x
XI4 net44 sync gnd vddp / inv_32x
XI2 ADCo BC Co Cob D<11> D<10> D<9> D<8> D<7> D<6> D<5> D<4> D<3> D<2> D<1> 
+ D<0> Ho PO<11> PO<10> PO<9> PO<8> PO<7> PO<6> PO<5> PO<4> PO<3> PO<2> PO<1> 
+ PO<0> RN Sa ck gnd lat vdd1p2 vddp / sarlogic2
XI0 gnd ib am ap lat Cob on Co vdda1p2 / comp2
.ENDS

